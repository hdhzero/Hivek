library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.hivek_pack.all;

entity hivek is
    port (
        clock : in std_logic;
        reset : in std_logic
    );
end hivek;

architecture hivek_arch of hivek is
begin
end hivek_arch;
