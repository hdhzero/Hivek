library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ikev is
    port (
        clock : in std_logic;
        reset : in std_logic
    );
end ikev;

architecture ikev_arch of ikev is
begin
end ikev_arch;
